proccess(clk)
begin
  case STATE is
    when s0 =>
      a = '1';
  end case;
end proccess;
